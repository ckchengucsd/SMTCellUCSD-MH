* CDL netlist for PROBE3.0
* Author: Minsoo Kim
* Based on ASAP7 CDL netlist
* 41 cell masters
* AND2_{X1,X2}, AND3_{X1,X2}, AOI21_{X1,X2}, AOI22_{X1,X2}, BUF_{X1,X2,X4,X8}, DFFHQN_X1, DFFRNQ_X1, LHQ_X1,
* INV_{X1,X2,X4,X8}, MUX2_X1, NAND2_{X1,X2}, NAND3_{X1,X2}, NAND4_{X1,X2}, NOR2_{X1,X2}, 
* NOR3_{X1,X2}, NOR4_{X1,X2}, OAI21_{X1,X2}, OAI22_{X1,X2}, OR2_{X1,X2}, OR3_{X1,X2}, XOR2_X1

* DGSB

.SUBCKT AND2_X1 A1 A2 VDD VSS Z
MM4 Z net10 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net10 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 net10 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 Z net10 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 net20 A2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net10 A1 net20 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AND2_X2 A1 A2 VDD VSS Z
MM4 Z net10 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 net10 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 Z net10 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net20 A2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net10 A1 net20 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS   

.SUBCKT AND2_X2Tr8 A1 A2 VDD VSS Z
*.PININFO
MM4 Z net10 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 net10 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 Z net10 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net20 A2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net10 A1 net20 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AND3_X1 A1 A2 A3 VDD VSS Z
MM7 Z net10 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 net10 A3 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net10 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net10 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 Z net10 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net30 A3 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net20 A2 net30 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net10 A1 net20 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AND3_X2 A1 A2 A3 VDD VSS Z
MM7 Z net10 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 net10 A3 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net10 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net10 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 Z net10 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 net30 A3 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net20 A2 net30 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net10 A1 net20 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AND3_X2Tr10 A1 A2 A3 VDD VSS Z
MM7 Z net10 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 net10 A3 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net10 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net10 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 Z net10 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 net30 A3 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net20 A2 net30 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net10 A1 net20 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AOI21_X1 A1 A2 B VDD VSS ZN
MM5 ZN B VSS VSS nmos_rvt w=23.00n l=16n nfin=1
MM4 net2 A1 ZN VSS nmos_rvt w=23.00n l=16n nfin=1
MM3 net2 A2 VSS VSS nmos_rvt w=23.00n l=16n nfin=1
MM2 net6 B VDD VDD pmos_rvt w=23.00n l=16n nfin=1
MM1 net6 A1 ZN VDD pmos_rvt w=23.00n l=16n nfin=1
MM0 net6 A2 ZN VDD pmos_rvt w=23.00n l=16n nfin=1
.ENDS

.SUBCKT AOI21_X2Tr12 A1 A2 B VDD VSS ZN
MM5 VSS B ZN VSS nmos_rvt w=46.00n l=16n nfin=2
MM4 ZN A1 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM3 VSS A2 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM2 VDD B net6 VDD pmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A1 net6 VDD pmos_rvt w=46.00n l=16n nfin=2
MM0 ZN A2 net6 VDD pmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT AOI21_X2 A1 A2 B VDD VSS ZN
MM5 VSS B ZN VSS nmos_rvt w=46.00n l=16n nfin=2
MM4 ZN A1 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM3 VSS A2 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM2 VDD B net6 VDD pmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A1 net6 VDD pmos_rvt w=46.00n l=16n nfin=2
MM0 ZN A2 net6 VDD pmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT AOI22_X1 A1 A2 B1 B2 VDD VSS ZN
MM7 net1 B2 VSS VSS nmos_rvt w=46.00n l=16n nfin=2
MM6 ZN B1 net1 VSS nmos_rvt w=46.00n l=16n nfin=2
MM5 net0 A1 ZN VSS nmos_rvt w=46.00n l=16n nfin=2
MM4 VSS A2 net0 VSS nmos_rvt w=46.00n l=16n nfin=2
MM3 net2 B2 VDD VDD pmos_rvt w=46.00n l=16n nfin=2
MM2 VDD B1 net2 VDD pmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A1 net2 VDD pmos_rvt w=46.00n l=16n nfin=2
MM0 net2 A2 ZN VDD pmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT AOI22_X2 A1 A2 B1 B2 VDD VSS ZN
MM7 net1 B2 VSS VSS nmos_rvt w=92.00n l=16n nfin=4
MM6 ZN B1 net1 VSS nmos_rvt w=92.00n l=16n nfin=4
MM5 net0 A1 ZN VSS nmos_rvt w=92.00n l=16n nfin=4
MM4 VSS A2 net0 VSS nmos_rvt w=92.00n l=16n nfin=4
MM3 net2 B2 VDD VDD pmos_rvt w=92.00n l=16n nfin=4
MM2 VDD B1 net2 VDD pmos_rvt w=92.00n l=16n nfin=4
MM1 ZN A1 net2 VDD pmos_rvt w=92.00n l=16n nfin=4
MM0 net2 A2 ZN VDD pmos_rvt w=92.00n l=16n nfin=4
.ENDS

.SUBCKT AOI22_X2Tr16 A1 A2 B1 B2 VDD VSS ZN
MM7 net1 B2 VSS VSS nmos_rvt w=46.00n l=16n nfin=2
MM6 ZN B1 net1 VSS nmos_rvt w=46.00n l=16n nfin=2
MM5 net0 A1 ZN VSS nmos_rvt w=46.00n l=16n nfin=2
MM4 VSS A2 net0 VSS nmos_rvt w=46.00n l=16n nfin=2
MM3 net2 B2 VDD VDD pmos_rvt w=46.00n l=16n nfin=2
MM2 VDD B1 net2 VDD pmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A1 net2 VDD pmos_rvt w=46.00n l=16n nfin=2
MM0 net2 A2 ZN VDD pmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT BUF_X1 I VDD VSS Z
MM3 Z IN VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 IN I VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 Z IN VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 IN I VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT BUF_X2 I VDD VSS Z
MM3 Z IN VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 IN I VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 Z IN VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 IN I VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT BUF_X4 I VDD VSS Z
MM3 Z IN VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM2 IN I VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM0 Z IN VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM1 IN I VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT BUF_X4Tr6 I VDD VSS Z
MM3 Z IN VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM2 IN I VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM0 Z IN VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM1 IN I VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT BUF_X8 I VDD VSS Z
MM3 Z IN VSS VSS nmos_rvt w=184.0n l=16n nfin=8
MM2 IN I VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM0 Z IN VDD VDD pmos_rvt w=184.0n l=16n nfin=8
MM1 IN I VDD VDD pmos_rvt w=92.0n l=16n nfin=4
.ENDS

.SUBCKT BUF_X8Tr6 I VDD VSS Z
MM3 Z IN VSS VSS nmos_rvt w=184.0n l=16n nfin=8
MM2 IN I VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM0 Z IN VDD VDD pmos_rvt w=184.0n l=16n nfin=8
MM1 IN I VDD VDD pmos_rvt w=92.0n l=16n nfin=4
.ENDS

.SUBCKT DFFHQN_X1 CLK D VDD VSS QN
MM4 net10 net3 net12 VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 VSS D net12 VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 VSS net10 net8 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 VSS net8 net9 VSS nmos_rvt w=23.0n l=16n nfin=1
MM9 net10 net4 net9 VSS nmos_rvt w=23.0n l=16n nfin=1
MM12 net8 net4 net1 VSS nmos_rvt w=23.0n l=16n nfin=1
MM14 net7 net1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM16 VSS net7 net6 VSS nmos_rvt w=23.0n l=16n nfin=1
MM17 net1 net3 net6 VSS nmos_rvt w=23.0n l=16n nfin=1
MM20 net3 CLK VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM23 net4 net3 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM24 QN net1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 VDD D net16 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net10 net4 net16 VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 VDD net10 net8 VDD pmos_rvt w=23.0n l=16n nfin=1
MM10 net10 net3 net15 VDD pmos_rvt w=23.0n l=16n nfin=1
MM11 VDD net8 net15 VDD pmos_rvt w=23.0n l=16n nfin=1
MM13 net8 net3 net1 VDD pmos_rvt w=23.0n l=16n nfin=1
MM15 net7 net1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM18 net1 net4 net14 VDD pmos_rvt w=23.0n l=16n nfin=1
MM19 VDD net7 net14 VDD pmos_rvt w=23.0n l=16n nfin=1
MM21 net3 CLK VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM22 net4 net3 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM25 QN net1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT DFFHQNEQFIN_X1 CLK D VDD VSS QN
MM4 net10 net3 net12 VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 VSS D net12 VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 VSS net10 net8 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 VSS net8 net9 VSS nmos_rvt w=23.0n l=16n nfin=1
MM9 net10 net4 net9 VSS nmos_rvt w=23.0n l=16n nfin=1
MM12 net8 net4 net1 VSS nmos_rvt w=23.0n l=16n nfin=1
MM14 net7 net1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM16 VSS net7 net6 VSS nmos_rvt w=23.0n l=16n nfin=1
MM17 net1 net3 net6 VSS nmos_rvt w=23.0n l=16n nfin=1
MM20 net3 CLK VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM23 net4 net3 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM24 QN net1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 VDD D net16 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net10 net4 net16 VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 VDD net10 net8 VDD pmos_rvt w=23.0n l=16n nfin=1
MM10 net10 net3 net15 VDD pmos_rvt w=23.0n l=16n nfin=1
MM11 VDD net8 net15 VDD pmos_rvt w=23.0n l=16n nfin=1
MM13 net8 net3 net1 VDD pmos_rvt w=23.0n l=16n nfin=1
MM15 net7 net1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM18 net1 net4 net14 VDD pmos_rvt w=23.0n l=16n nfin=1
MM19 VDD net7 net14 VDD pmos_rvt w=23.0n l=16n nfin=1
MM21 net3 CLK VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM22 net4 net3 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM25 QN net1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT INV_X1 I VDD VSS ZN
MM0 ZN I VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 ZN I VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS


.SUBCKT INV_X2 I VDD VSS ZN
MM0 ZN I VSS VSS nmos_rvt w=92.00n l=16n nfin=4
MM1 ZN I VDD VDD pmos_rvt w=92.00n l=16n nfin=4
.ENDS

.SUBCKT INV_X4 I VDD VSS ZN
MM0 ZN I VSS VSS nmos_rvt w=92.00n l=16n nfin=4
MM1 ZN I VDD VDD pmos_rvt w=92.00n l=16n nfin=4
.ENDS

.SUBCKT INV_X8 I VDD VSS ZN
MM0 ZN I VSS VSS nmos_rvt w=184.0n l=16n nfin=8
MM1 ZN I VDD VDD pmos_rvt w=184.00n l=16n nfin=8
.ENDS


.SUBCKT MUX2_X1 I0 I1 S VDD VSS Z
MM11 Z net5 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM10 VSS I0 net6 VSS nmos_rvt w=23.0n l=16n nfin=1
MM9 net6 net2 net5 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 net5 S net4 VSS nmos_rvt w=23.0n l=16n nfin=1
MM7 VSS I1 net4 VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 net2 S VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 Z net5 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 VDD I0 net11 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 net11 S net5 VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net5 net2 net10 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 VDD I1 net10 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 net2 S VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS


.SUBCKT NAND2_X1 A1 A2 VDD VSS ZN
MM3 net16 A2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 ZN A1 net16 VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 ZN A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 ZN A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT NAND2_X2 A1 A2 VDD VSS ZN
MM3 net16 A2 VSS VSS nmos_rvt w=92.00n l=16n nfin=4
MM2 ZN A1 net16 VSS nmos_rvt w=92.00n l=16n nfin=4
MM1 ZN A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 ZN A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NAND2_X2Tr8 A1 A2 VDD VSS ZN
MM3 net16 A2 VSS VSS nmos_rvt w=46.00n l=16n nfin=2
MM2 ZN A1 net16 VSS nmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 ZN A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NAND3_X1 A1 A2 A3 VDD VSS ZN
MM5 net17 A3 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 net16 A2 net17 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 ZN A1 net16 VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 ZN A3 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 ZN A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 ZN A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT NAND3_X2 A1 A2 A3 VDD VSS ZN
MM5 net17 A3 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 net16 A2 net17 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 ZN A1 net16 VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 ZN A3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 ZN A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 ZN A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NAND3_X2Tr12 A1 A2 A3 VDD VSS ZN
MM5 net17 A3 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 net16 A2 net17 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 ZN A1 net16 VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 ZN A3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 ZN A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 ZN A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NAND4_X1 A1 A2 A3 A4 VDD VSS ZN
MM7 net18 A4 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 net17 A3 net18 VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 net16 A2 net17 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 ZN A1 net16 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 ZN A4 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 ZN A3 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 ZN A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 ZN A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT NAND4_X2 A1 A2 A3 A4 VDD VSS ZN
MM7 net18 A4 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 net17 A3 net18 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 net16 A2 net17 VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 ZN A1 net16 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 ZN A4 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 ZN A3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 ZN A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 ZN A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NAND4_X2Tr16 A1 A2 A3 A4 VDD VSS ZN
MM7 net18 A4 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 net17 A3 net18 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 net16 A2 net17 VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 ZN A1 net16 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 ZN A4 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 ZN A3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 ZN A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 ZN A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NOR2_X1 A1 A2 VDD VSS ZN
MM3 VSS A1 ZN VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 VSS A2 ZN VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net16 A1 ZN VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A2 net16 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT NOR2_X2 A1 A2 VDD VSS ZN
MM3 VSS A1 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 VSS A2 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM1 net16 A1 ZN VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A2 net16 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NOR2_X2Tr8 A1 A2 VDD VSS ZN
MM3 VSS A1 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 VSS A2 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM1 net16 A1 ZN VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A2 net16 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NOR3_X1 A1 A2 A3 VDD VSS ZN
MM5 VSS A1 ZN VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 VSS A2 ZN VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 VSS A3 ZN VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net20 A1 ZN VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net10 A2 net20 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A3 net10 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT NOR3_X2 A1 A2 A3 VDD VSS ZN
MM5 VSS A1 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A2 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 VSS A3 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 net20 A1 ZN VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 A2 net20 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A3 net10 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NOR3_X2Tr12 A1 A2 A3 VDD VSS ZN
MM5 VSS A1 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A2 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 VSS A3 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 net20 A1 ZN VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 A2 net20 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A3 net10 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NOR4_X1 A1 A2 A3 A4 VDD VSS ZN
MM7 VSS A1 ZN VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 VSS A2 ZN VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 VSS A3 ZN VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 VSS A4 ZN VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 net30 A1 ZN VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net20 A2 net30 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net10 A3 net20 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A4 net10 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT NOR4_X2 A1 A2 A3 A4 VDD VSS ZN
MM7 VSS A1 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS A2 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 VSS A3 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A4 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net30 A1 ZN VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net20 A2 net30 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 A3 net20 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A4 net10 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NOR4_X2Tr16 A1 A2 A3 A4 VDD VSS ZN
MM7 VSS A1 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS A2 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 VSS A3 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A4 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net30 A1 ZN VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net20 A2 net30 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 A3 net20 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A4 net10 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT OAI21_X1 A1 A2 B VDD VSS ZN
MM5 VDD B ZN VDD pmos_rvt w=23.00n l=16n nfin=1
MM3 ZN A1 net7 VDD pmos_rvt w=23.00n l=16n nfin=1
MM4 VDD A2 net7 VDD pmos_rvt w=23.00n l=16n nfin=1
MM2 VSS B net0 VSS nmos_rvt w=23.00n l=16n nfin=1
MM0 ZN A1 net0 VSS nmos_rvt w=23.00n l=16n nfin=1
MM1 ZN A2 net0 VSS nmos_rvt w=23.00n l=16n nfin=1
.ENDS

.SUBCKT OAI21_X2 A1 A2 B VDD VSS ZN
MM5 VDD B ZN VDD pmos_rvt w=46.00n l=16n nfin=2
MM3 ZN A1 net7 VDD pmos_rvt w=46.00n l=16n nfin=2
MM4 VDD A2 net7 VDD pmos_rvt w=46.00n l=16n nfin=2
MM2 VSS B net0 VSS nmos_rvt w=46.00n l=16n nfin=2
MM0 ZN A1 net0 VSS nmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A2 net0 VSS nmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT OAI21_X2Tr12 A1 A2 B VDD VSS ZN
MM5 VDD B ZN VDD pmos_rvt w=46.00n l=16n nfin=2
MM3 ZN A1 net7 VDD pmos_rvt w=46.00n l=16n nfin=2
MM4 VDD A2 net7 VDD pmos_rvt w=46.00n l=16n nfin=2
MM2 VSS B net0 VSS nmos_rvt w=46.00n l=16n nfin=2
MM0 ZN A1 net0 VSS nmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A2 net0 VSS nmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT OAI22_X1 A1 A2 B1 B2 VDD VSS ZN
MM7 VDD B2 net8 VDD pmos_rvt w=46.00n l=16n nfin=2
MM6 ZN B1 net8 VDD pmos_rvt w=46.00n l=16n nfin=2
MM4 net9 A1 ZN VDD pmos_rvt w=46.00n l=16n nfin=2
MM5 VDD A2 net9 VDD pmos_rvt w=46.00n l=16n nfin=2
MM3 VSS B2 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM2 VSS B1 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM0 ZN A1 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A2 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT OAI22_X2 A1 A2 B1 B2 VDD VSS ZN
MM7 VDD B2 net8 VDD pmos_rvt w=92.00n l=16n nfin=4
MM6 ZN B1 net8 VDD pmos_rvt w=92.00n l=16n nfin=4
MM4 net9 A1 ZN VDD pmos_rvt w=92.00n l=16n nfin=4
MM5 VDD A2 net9 VDD pmos_rvt w=92.00n l=16n nfin=4
MM3 VSS B2 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
MM2 VSS B1 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
MM0 ZN A1 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
MM1 ZN A2 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
.ENDS

.SUBCKT OAI22_X2Tr16 A1 A2 B1 B2 VDD VSS ZN
MM7 VDD B2 net8 VDD pmos_rvt w=46.00n l=16n nfin=2
MM6 ZN B1 net8 VDD pmos_rvt w=46.00n l=16n nfin=2
MM4 net9 A1 ZN VDD pmos_rvt w=46.00n l=16n nfin=2
MM5 VDD A2 net9 VDD pmos_rvt w=46.00n l=16n nfin=2
MM3 VSS B2 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM2 VSS B1 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM0 ZN A1 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A2 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT OR2_X1 A1 A2 VDD VSS Z
MM5 Z net2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 VSS A1 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 VSS A2 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 Z net2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net2 A1 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A2 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OR2_X2 A1 A2 VDD VSS Z
MM5 Z net2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A1 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 VSS A2 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 Z net2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net2 A1 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A2 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OR2_X2Tr8 A1 A2 VDD VSS Z
MM5 Z net2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A1 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 VSS A2 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 Z net2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net2 A1 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A2 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OR3_X1 A1 A2 A3 VDD VSS Z
MM7 Z net2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 VSS A1 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 VSS A2 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 VSS A3 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 Z net2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net2 A1 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net7 A2 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A3 net7 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OR3_X2 A1 A2 A3 VDD VSS Z
MM7 Z net2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS A1 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 VSS A2 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 VSS A3 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 Z net2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net2 A1 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net7 A2 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A3 net7 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OR3_X2Tr10 A1 A2 A3 VDD VSS Z
MM7 Z net2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS A1 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 VSS A2 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 VSS A3 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 Z net2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net2 A1 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net7 A2 net6 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A3 net7 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT XOR2_X1 A1 A2 VDD VSS Z
MM9 VSS A2 net5 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 net5 A1 Z VSS nmos_rvt w=23.0n l=16n nfin=1
MM7 VSS net2 Z VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 VSS A1 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 VSS A2 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 Z A2 net8 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 Z A1 net8 VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 VDD net2 net8 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net2 A1 net7 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD A2 net7 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS


.SUBCKT DFFRNQ_X1 D RN CK Q VDD VSS 
MM27 VSS CK ncki VSS nmos_rvt w=23.0n l=16n nfin=1
MM26 cki ncki VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM25 net10 D VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM24 net1 ncki net10 VSS nmos_rvt w=23.0n l=16n nfin=1
MM23 net15 cki net1 VSS nmos_rvt w=23.0n l=16n nfin=1
MM22 net12 net2 net15 VSS nmos_rvt w=23.0n l=16n nfin=1
MM21 VSS RN net12 VSS nmos_rvt w=23.0n l=16n nfin=1
MM20 net2 net1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM19 net8 cki net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM18 net11 ncki net8 VSS nmos_rvt w=23.0n l=16n nfin=1
MM17 VSS net4 net11 VSS nmos_rvt w=23.0n l=16n nfin=1
MM16 net0 RN VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM15 net4 net8 net0 VSS nmos_rvt w=23.0n l=16n nfin=1
MM14 VSS net4 Q VSS nmos_rvt w=23.0n l=16n nfin=1
MM13 VDD CK ncki VDD pmos_rvt w=23.0n l=16n nfin=1
MM12 cki ncki VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM11 net10 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM10 net1 cki net10 VDD pmos_rvt w=23.0n l=16n nfin=1
MM9 net9 ncki net1 VDD pmos_rvt w=23.0n l=16n nfin=1
MM8 VDD net2 net9 VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 net9 RN VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 net2 net1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net8 ncki net2 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net11 cki net8 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 VDD net4 net11 VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net4 RN VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 VDD net8 net4 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD net4 Q VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS 

.SUBCKT DFFRNQEQFIN_X1 D RN CK Q VDD VSS 
MM27 VSS CK ncki VSS nmos_rvt w=23.0n l=16n nfin=1
MM26 cki ncki VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM25 net10 D VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM24 net1 ncki net10 VSS nmos_rvt w=23.0n l=16n nfin=1
MM23 net15 cki net1 VSS nmos_rvt w=23.0n l=16n nfin=1
MM22 net12 net2 net15 VSS nmos_rvt w=23.0n l=16n nfin=1
MM21 VSS RN net12 VSS nmos_rvt w=23.0n l=16n nfin=1
MM20 net2 net1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM19 net8 cki net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM18 net11 ncki net8 VSS nmos_rvt w=23.0n l=16n nfin=1
MM17 VSS net4 net11 VSS nmos_rvt w=23.0n l=16n nfin=1
MM16 net0 RN VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM15 net4 net8 net0 VSS nmos_rvt w=23.0n l=16n nfin=1
MM14 VSS net4 Q VSS nmos_rvt w=23.0n l=16n nfin=1
MM13 VDD CK ncki VDD pmos_rvt w=23.0n l=16n nfin=1
MM12 cki ncki VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM11 net10 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM10 net1 cki net10 VDD pmos_rvt w=23.0n l=16n nfin=1
MM9 net9 ncki net1 VDD pmos_rvt w=23.0n l=16n nfin=1
MM8 VDD net2 net9 VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 net9 RN VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 net2 net1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net8 ncki net2 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net11 cki net8 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 VDD net4 net11 VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net4 RN VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 VDD net8 net4 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD net4 Q VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS 

.SUBCKT LHQ_X1 D E Q VDD VSS 
MM15 net4 E VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM14 net7 net4 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM13 net3 D VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM12 net5 net7 net3 VSS nmos_rvt w=23.0n l=16n nfin=1
MM11 net2 net4 net5 VSS nmos_rvt w=23.0n l=16n nfin=1
MM10 VSS net6 net2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM9 net6 net5 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 Q net5 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM7 net4 E VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 net7 net4 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net1 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net5 net4 net1 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 net0 net7 net5 VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 VDD net6 net0 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net6 net5 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 Q net5 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS 

.SUBCKT A2O1A1O1I_X1 A1 A2 B C D VDD VSS Y
MM5 net4 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM8 net15 C VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 net4 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM9 Y D net15 VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 net15 B net4 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 Y D VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net25 A2 net12 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 Y B net12 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 Y A1 net25 VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net12 C VSS VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT A2O1A1I_X1 A1 A2 B C VDD VSS Y
MM7 net06 B VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 Y C net06 VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net015 A2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net06 A1 net015 VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 Y C VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 Y B net2 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net2 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 net2 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AND4_X1 A B C D VDD VSS Y
MM8 Y net12 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 net12 A VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 net12 B VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net12 C VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net12 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM9 Y net12 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 pd3 A VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 pd2 B pd3 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 pd1 C pd2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net12 D pd1 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AND4_X2 A B C D VDD VSS Y
MM8 Y net12 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM7 net12 A pd1 VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 pd1 B pd2 VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 pd2 C pd3 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 pd3 D VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM9 Y net12 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM3 net12 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net12 C VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net12 B VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 net12 A VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AND5_X1 A B C D E VDD VSS Y
MM11 Y net011 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 net29 E VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 net30 D net29 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 net024 B net023 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net011 A net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 net023 C net30 VSS nmos_rvt w=23.0n l=16n nfin=1
MM9 net011 E VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM8 net011 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 net011 C VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net011 B VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 Y net011 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM10 net011 A VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AND5_X2 A B C D E VDD VSS Y
MM11 VSS net024 Y VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS E net027 VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 net027 D net29 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 net30 B net023 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net023 A net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 net29 C net30 VSS nmos_rvt w=23.0n l=16n nfin=1
MM9 VDD E net024 VDD pmos_rvt w=23.0n l=16n nfin=1
MM8 VDD D net024 VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 VDD C net024 VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 VDD B net024 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 VDD net024 Y VDD pmos_rvt w=46.0n l=16n nfin=2
MM10 VDD A net024 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OR4_X1 A B C D VDD VSS Y
MM9 Y net12 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 net12 D VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net12 C VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net12 B VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net12 A VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 Y net12 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 net12 A pd1 VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 pd1 B pd2 VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 pd2 C pd3 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 pd3 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OR4_X2 A B C D VDD VSS Y
MM9 Y net12 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net12 D VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net12 C VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net12 B VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net12 A VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 Y net12 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM7 net12 A pd1 VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 pd1 B pd2 VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 pd2 C pd3 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 pd3 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OR5_X1 A B C D E VDD VSS Y
MM9 VSS E net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 VSS D net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM7 VSS C net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 VSS B net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 VSS net024 Y VSS nmos_rvt w=23.0n l=16n nfin=1
MM10 VSS A net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM11 VDD net024 Y VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 VDD E net027 VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net027 D net29 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net30 B net023 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 net023 A net024 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 net29 C net30 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OR5_X2 A B C D E VDD VSS Y
MM9 VSS E net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 VSS D net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM7 VSS C net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 VSS B net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 VSS net024 Y VSS nmos_rvt w=46.0n l=16n nfin=2
MM10 VSS A net024 VSS nmos_rvt w=23.0n l=16n nfin=1
MM11 VDD net024 Y VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 VDD E net027 VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net027 D net29 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net30 B net023 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 net023 A net024 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 net29 C net30 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AO21_X1 A1 A2 B VDD VSS Y
MM7 Y net16 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 net16 B VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 net16 A1 net29 VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net29 A2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 Y net16 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net18 A2 net16 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD B net18 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net18 A1 net16 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AO21_X2 A1 A2 B VDD VSS Y
MM7 Y net16 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 net16 B VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 net16 A1 net29 VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net29 A2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 Y net16 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM5 net18 A2 net16 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 VDD B net18 VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net18 A1 net16 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AO22_X1 A1 A2 B1 B2 VDD VSS Y
MM5 net18 B2 net13 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net18 B1 net13 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 net13 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 Y net18 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net13 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM9 net29 B1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 net30 A1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM7 net18 B2 net29 VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 net18 A2 net30 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 Y net18 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT AO22_X2 A1 A2 B1 B2 VDD VSS Y
MM5 net18 B2 net13 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net18 B1 net13 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 net13 A2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 Y net18 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net13 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM9 net29 B1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 net30 A1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM7 net18 B2 net29 VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 net18 A2 net30 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 Y net18 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT DLL_X1 CLK D Q VDD VSS
MM23 clkb clkn VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 pd1 D VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 MH clkn pd1 VSS nmos_rvt w=23.0n l=16n nfin=1
MM20 clkn CLK VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM24 Q MH VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 net085 MH VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM9 MH clkb pd3 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 pd3 net085 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM22 clkb clkn VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 MH clkb pu1 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 pu1 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM25 Q MH VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM21 clkn CLK VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 net085 MH VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM11 pd2 net085 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM10 MH clkn pd2 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT DLL_X2 CLK D Q VDD VSS
MM23 clkb clkn VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 pd1 D VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 MH clkn pd1 VSS nmos_rvt w=23.0n l=16n nfin=1
MM24 Q MH VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM20 clkn CLK VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 net085 MH VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM9 MH clkb pd3 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 pd3 net085 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM11 pd2 net085 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM10 MH clkn pd2 VDD pmos_rvt w=23.0n l=16n nfin=1
MM22 clkb clkn VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 MH clkb pu1 VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 pu1 D VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM21 clkn CLK VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM25 Q MH VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM7 net085 MH VDD VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT O2A1O1I_X1 A1 A2 B C VDD VSS Y
MM7 net010 B VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 Y C net010 VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 net010 A2 net019 VDD pmos_rvt w=23.0n l=16n nfin=1
MM4 net019 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM3 Y C VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net022 B VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 Y A2 net022 VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 Y A1 net022 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OA21_X1 A1 A2 B VDD VSS Y
MM3 Y net25 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net25 B VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net25 A2 net27 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 net27 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 Y net25 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 net11 B VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 net25 A2 net11 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 net25 A1 net11 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OA21_X2 A1 A2 B VDD VSS Y
MM3 Y net25 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net25 B VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM1 net25 A2 net27 VDD pmos_rvt w=23.0n l=16n nfin=1
MM0 net27 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 Y net25 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 net11 B VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 net25 A2 net11 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 net25 A1 net11 VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OA22_X1 A1 A2 B1 B2 VDD VSS Y
MM9 Y net033 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 net3 B2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net033 A2 net3 VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net3 B1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net033 A1 net3 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 net13 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM11 net033 A2 net13 VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 net14 B1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 Y net033 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM10 net033 B2 net14 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT OA22_X2 A1 A2 B1 B2 VDD VSS Y
MM9 Y net033 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net3 B2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM2 net033 A2 net3 VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net3 B1 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 net033 A1 net3 VSS nmos_rvt w=23.0n l=16n nfin=1
MM8 net13 A1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM11 net033 A2 net13 VDD pmos_rvt w=23.0n l=16n nfin=1
MM6 net14 B1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM5 Y net033 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM10 net033 B2 net14 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT TIELO_X1 L VDD VSS
MM1 net9 L VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 L net9 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT TIELO_X2 L VDD VSS
MM1 net9 L VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 L net9 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT TIEHI_X1 H VDD VSS
MM1 H net7 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM2 net7 H VSS VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS

.SUBCKT TIEHI_X2 H VDD VSS
MM1 H net7 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net7 H VSS VSS nmos_rvt w=23.0n l=16n nfin=1
.ENDS


.SUBCKT AOI2222_Xp33 A1 A2 B1 B2 C1 C2 D1 D2 VDD VSS Y
MM14 net48 D2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM13 Y D1 net48 VSS nmos_rvt w=23.0n l=16n nfin=1
MM6 net50 C2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM5 Y C1 net50 VSS nmos_rvt w=23.0n l=16n nfin=1
MM4 net51 B2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM3 Y B1 net51 VSS nmos_rvt w=23.0n l=16n nfin=1
MM1 net49 A2 VSS VSS nmos_rvt w=23.0n l=16n nfin=1
MM0 Y A1 net49 VSS nmos_rvt w=23.0n l=16n nfin=1
MM16 net11 D2 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM15 net11 D1 VDD VDD pmos_rvt w=23.0n l=16n nfin=1
MM12 Y A2 net53 VDD pmos_rvt w=23.0n l=16n nfin=1
MM11 net53 B2 net27 VDD pmos_rvt w=23.0n l=16n nfin=1
MM10 net27 C2 net11 VDD pmos_rvt w=23.0n l=16n nfin=1
MM9 Y A1 net53 VDD pmos_rvt w=23.0n l=16n nfin=1
MM8 net53 B1 net27 VDD pmos_rvt w=23.0n l=16n nfin=1
MM7 net27 C1 net11 VDD pmos_rvt w=23.0n l=16n nfin=1
.ENDS
