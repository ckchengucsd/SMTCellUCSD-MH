VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;

SITE coresite
    SIZE 0.0450 BY -0.0240 ;
    CLASS CORE ;
    SYMMETRY Y ;
END coresite

MACRO BUF_X4Tr6_5T_2F_45CPP_24M0P_30M1P_24M2P_2MPO_ET_BPR
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X4Tr6_5T_2F_45CPP_24M0P_30M1P_24M2P_2MPO_ET_BPR 0 0 ;
  SIZE 0.1800 BY 0.2400 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0225 0.1080 0.0375 0.0360 ;
    END
  END Z
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1125 0.1320 0.1275 0.0840 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.2330 0.1800 0.2470 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0070 0.1800 0.0070 ;
    END
  END VSS
  OBS
      LAYER M1 ;
        RECT 0.0525 0.1320 0.0675 0.0600 ;
  END
END BUF_X4Tr6_5T_2F_45CPP_24M0P_30M1P_24M2P_2MPO_ET_BPR

END LIBRARY
